//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab8(input               CLOCK_50,
            input        [3:0]  KEY,          //bit 0 is set up as Reset
            input logic  [3:0]  SW,
            output logic [6:0]  HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7,

            // VGA Interface 
            output logic [7:0]  VGA_R,        //VGA Red
                                VGA_G,        //VGA Green
                                VGA_B,        //VGA Blue
            output logic        VGA_CLK,      //VGA Clock
                                VGA_SYNC_N,   //VGA Sync signal
                                VGA_BLANK_N,  //VGA Blank signal
                                VGA_VS,       //VGA virtical sync signal
                                VGA_HS,       //VGA horizontal sync signal

            // CY7C67200 Interface
            inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
            output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
            output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                OTG_RD_N,     //CY7C67200 Write
                                OTG_WR_N,     //CY7C67200 Read
                                OTG_RST_N,    //CY7C67200 Reset
            input               OTG_INT,      //CY7C67200 Interrupt

            // SDRAM Interface for Nios II Software
            output logic [12:0]  DRAM_ADDR,    //SDRAM Address 13 Bits
            inout  wire  [31:0]  DRAM_DQ,      //SDRAM Data 32 Bits
            output logic [1:0]   DRAM_BA,      //SDRAM Bank Address 2 Bits
            output logic [3:0]   DRAM_DQM,     //SDRAM Data Mast 4 Bits
            output logic         DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK,     //SDRAM Clock

            input logic         AUD_ADCDAT,
            input logic         AUD_BCLK,
            input logic         AUD_ADCLRCK,
            input logic         AUD_DACLRCK,
            output logic        AUD_DACDAT,
            output logic        AUD_XCK,
            output logic        I2C_SCLK,
            output logic        I2C_SDAT,

            output logic            FL_WE_N,   //FLASH Write Enable
                                    FL_RST_N,  //FLASH Reset
                                    FL_WP_N,   //FLASH Write Protect
                                    FL_CE_N,   //FLASH Chip Enable
                                    FL_OE_N,   //FLASH Output Enable
            input  logic            FL_RY,     //FLASH Ready Busy Output
            output logic  [22:0]    FL_ADDR,   //FLASH Address
            input  logic  [7 :0]    FL_DQ      //FLASH Data

                    );
    
    logic Reset_h, Clk;
    logic [15:0] keycode;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs;
     
     logic [9:0] World_X, World_Y;
     logic is_sprite;
     
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),    
                            .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     lab8_soc nios_system(
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w)
    );
  
    // Use PLL to generate the 25MHZ VGA_CLK. Do not modify it.
    // vga_clk vga_clk_instance(
    //     .clk_clk(Clk),
    //     .reset_reset_n(1'b1),
    //     .altpll_0_c0_clk(VGA_CLK),
    //     .altpll_0_areset_conduit_export(),    
    //     .altpll_0_locked_conduit_export(),
    //     .altpll_0_phasedone_conduit_export()
    // );
    always_ff @ (posedge Clk) begin
        if(Reset_h)
            VGA_CLK <= 1'b0;
        else
            VGA_CLK <= ~VGA_CLK;
    end
    
    audio audio_instance(.*);

    VGA_controller vga_controller_instance(.*,
                                                         .Reset(Reset_h),
                                                         .DrawX(World_X),
                                                         .DrawY(World_Y));
    
    sprite sprite_map(.*,
                              .is_sprite(is_sprite),
                              .Reset(Reset_h),
                              .frame_clk(VGA_VS),
                              .DrawX(World_X),
                              .DrawY(World_Y),
                              .Keycode(keycode[7:0]),
                              .run(SW[0])
                      );

    color_mapper color_instance(.*,
                                .Reset(Reset_h),
                                .run(SW[0]),
                                .DrawX(World_X),
                                .DrawY(World_Y));

	 // Display keycode on hex display
    HexDriver hex_inst_0 (keycode[3:0], HEX0);
    HexDriver hex_inst_1 (keycode[7:4], HEX1);
    // HexDriver hex0 (delay[3 :0 ], HEX0);
    // HexDriver hex1 (delay[7 :4 ], HEX1);
    // HexDriver hex2 (delay[11:8 ], HEX2);
    // HexDriver hex3 (delay[15:12], HEX3);
    // HexDriver hex4 (delay[19:16], HEX4);
    // HexDriver hex5 (delay[23:20], HEX5);
    // HexDriver hex6 (delay[27:24], HEX6);
    // HexDriver hex7 (delay[31:28], HEX7);
    
    /**************************************************************************************
        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
        Hidden Question #1/2:
        What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
             connect to the keyboard? List any two.  Give an answer in your Post-Lab.
    **************************************************************************************/
endmodule
